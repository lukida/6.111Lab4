library verilog;
use verilog.vl_types.all;
entity FSMTest is
end FSMTest;
