library verilog;
use verilog.vl_types.all;
entity FSMTest2 is
end FSMTest2;
