library verilog;
use verilog.vl_types.all;
entity FSMTest6 is
end FSMTest6;
