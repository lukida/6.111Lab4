library verilog;
use verilog.vl_types.all;
entity FSMTest3 is
end FSMTest3;
